* Sinusoidal voltage source

v1 a 0 sin(0 10 1MEG 0 0 0)
r1 a 0 1k
.tran 1n 2u
.plot tran v(a)
.end
